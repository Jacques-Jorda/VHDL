LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY multiplexer IS
	PORT (	E : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			C : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			S : OUT STD_LOGIC);
END ENTITY multiplexer;


ARCHITECTURE fdd_MPX OF multiplexer IS
BEGIN
	WITH C SELECT
		S <= 	E(0) WHEN "00",
				E(1) WHEN "01",
				E(2) WHEN "10",
				E(3) WHEN "11",
				'X' WHEN OTHERS;
END ARCHITECTURE fdd_MPX;
